package alu_types is
	type TYPE_OP is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, FUNCASL, FUNCASR, FUNCRL, FUNCRR);
end alu_types;